library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_128x17 is
    port (
        clk         : in std_logic;                 -- synchronous rom
        addr        : in unsigned(6 downto 0);      -- 128 addresses
        data_out    : out unsigned(16 downto 0)     -- 17 bits of data
    );
end entity;

architecture a_rom_128x17 of rom_128x17 is
    type mem is array (0 to 127) of unsigned(16 downto 0); -- 128 addresses, 17 bits of data
    constant rom_data: mem := (
        -- case addr => data
        0   => "1111" & "0000000000001",
        1   => "1111" & "0000000000100",
        2   => "0000" & "0000000000000",
        3   => "0000" & "0000000000000",
        4   => "0000" & "0000000000000",
        5   => "1111" & "0000000000111",
        6   => "0000" & "0000000000000",
        7   => "1111" & "0000000001010",
        8   => "0000" & "0000000000000",
        9   => "0000" & "0000000000000",
        10  => "1111" & "0000000000101",
        -- omitted cases
        others => (others => '0')
    );

begin
    process(clk)
    begin
        if(rising_edge(clk)) then
            data_out <= rom_data(to_integer(addr));
        end if;
    end process;
end architecture ;
