library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_128x17 is
    port (
        clk         : in std_logic;                 -- synchronous rom
        addr        : in unsigned(6 downto 0);      -- 128 addresses
        data_out    : out unsigned(16 downto 0)     -- 17 bits of data
    );
end entity;

architecture a_rom_128x17 of rom_128x17 is
    type mem is array (0 to 127) of unsigned(16 downto 0); -- 128 addresses, 17 bits of data
    constant rom_data: mem := (
        -- case addr => data
        0   => "0011" & "0000100001" & "001",               -- MOVEI.W #$33, D1         (0x06109)
        1   => "0011" & "0000000010" & "010",               -- MOVEI.W #$2, D2          (0x06012)
        2   => "0011" & "0000000001" & "011",               -- MOVEI.W #$1, D3          (0x0600B)

        3   => "1001" & "0000000" & "010" & "010",          -- loopX: MOVE.W D2, (D2)   (0x12012)
        4   => "0001" & "0000000" & "011" & "010",          -- ADD.W D3, D2             (0x0201A)
        5   => "0101" & "0000000" & "001" & "010",          -- CMP.W D1, D2             (0x0A00A)
        6   => "0111" & "00000"   & "0"   & "0000011",      -- BLT.S loopX              (0x0E003)

        7   => "0011" & "0000000100" & "010",               -- MOVEI.W #$4, D2          (0x06022)
        8   => "0011" & "0000000010" & "011",               -- MOVEI.W #$2, D3          (0x06013)
        9   => "1001" & "0000000" & "000" & "010",          -- loop2: MOVE.W D0, (D2)   (0x12002)
        10  => "0001" & "0000000" & "011" & "010",          -- ADD.W D3, D2             (0x0201A)
        11  => "0101" & "0000000" & "001" & "010",          -- CMP.W D1, D2             (0x0A00A)
        12  => "0111" & "00000"   & "0"   & "0001001",      -- BLT.S loop2              (0x0E009)

        13  => "0011" & "0000000110" & "010",               -- MOVEI.W #$6, D2          (0x06032)
        14  => "0011" & "0000000011" & "011",               -- MOVEI.W #$3, D3          (0x0601B)
        15  => "1001" & "0000000" & "000" & "010",          -- loop3: MOVE.W D0, (D2)   (0x12002)
        16  => "0001" & "0000000" & "011" & "010",          -- ADD.W D3, D2             (0x0201A)
        17  => "0101" & "0000000" & "001" & "010",          -- CMP.W D1, D2             (0x0A00A)
        18  => "0111" & "00000"   & "0"   & "0001111",      -- BLT.S loop3              (0x0E00F)

        19  => "0011" & "0000001010" & "010",               -- MOVEI.W #$10, D2         (0x06052)
        20  => "0011" & "0000000101" & "011",               -- MOVEI.W #$5, D3          (0x0602B)
        21  => "1001" & "0000000" & "000" & "010",          -- loop5: MOVE.W D0, (D2)   (0x12002)
        22  => "0001" & "0000000" & "011" & "010",          -- ADD.W D3, D2             (0x0201A)
        23  => "0101" & "0000000" & "001" & "010",          -- CMP.W D1, D2             (0x0A00A)
        24  => "0111" & "00000"   & "0"   & "0010101",      -- BLT.S loop5              (0x0E015)

        25  => "0011" & "0000100001" & "001",               -- MOVEI.W #$33, D1         (0x06109)
        26  => "0011" & "0000000010" & "010",               -- MOVEI.W #$2, D2          (0x06012)
        27  => "0011" & "0000000001" & "011",               -- MOVEI.W #$1, D3          (0x0600B)

        28  => "1000" & "0000000" & "010" & "100",          -- loopR: MOVE.W (D2), D4   (0x10014)
        29  => "0001" & "0000000" & "011" & "010",          -- ADD.W D3, D2             (0x0201A)
        30  => "0101" & "0000000" & "000" & "100",          -- CMP.W D0, D4             (0x0A004)
        31  => "0110" & "00000"   & "0"   & "0100010",      -- BEQ.S notPrime           (0x0C022)
        32  => "0100" & "0000000" & "100" & "101",          -- MOVE.W D4, D5            (0x08025)
        33  => "1111" & "00000"   & "0"   & "0011100",      -- JMP loopR                (0x1E01C)

        34  => "0101" & "0000000" & "010" & "001",          -- notPrime: CMP.W D2, D1   (0x0A011)
        35  => "0110" & "00000"   & "0"   & "1111111",      -- BEQ.S end                (0x0C07F)
        36  => "1111" & "00000"   & "0"   & "0011100",      -- JMP loopR                (0x1E01C)

        127 => "00000000000000000",                         -- end: NOP                 (0x00000)

        -- omitted cases
        others => (others => '0')
    );

begin
    process(clk)
    begin
        if(rising_edge(clk)) then
            data_out <= rom_data(to_integer(addr));
        end if;
    end process;
end architecture ;
