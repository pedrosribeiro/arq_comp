library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity processor is
    port (
        -- ports definition
    );
end entity;

architecture a_processor of processor is
    
begin
   
end architecture;